// Code your design here
module mux_2_1(
  input a,
  input b,
  input select,
  output y
);

  assign y = (select)?b:a;
endmodule