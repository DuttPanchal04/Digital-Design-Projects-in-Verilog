// Code your design here
// Code your design here
// Code your design here
// Code your design here
// Code your design here
module xor_gate(

	input a,
  	input b,
  	output y
  
);
  
  assign y = a^b;
  
endmodule